module main

fn main() {
	// files := walk_directory()

	// println(files)
	run()
}
