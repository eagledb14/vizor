module main




